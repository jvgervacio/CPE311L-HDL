primitive _2X1_MUX(
    output Y,
    input S, A, B
);
    table
      // S A B : Y
      0 0 ? : 0;
      0 1 ? : 1;
      1 ? 0 : 0;
      1 ? 1 : 1;
    endtable
endprimitive

module _8x1_MUX(
    output          Y,
    input [2:0]     S,
    input [7:0]     I
);
    wire [5:0] w;

    _2X1_MUX    
        mux0(w[0], S[0], I[0], I[1]),
        mux1(w[1], S[0], I[2], I[3]),
        mux2(w[2], S[0], I[4], I[5]),
        mux3(w[3], S[0], I[6], I[7]),

        mux4(w[4], S[1], w[0], w[1]),
        mux5(w[5], S[1], w[2], w[3]),

        mux6(   Y, S[2], w[4], w[5]);

endmodule

module exercise4_1;
    reg [7:0]   I;
    reg [2:0]   S;
    wire        Y;

    _8x1_MUX mux(Y, S, I);

    initial begin
            $display("8x1 MULTIPLEXER");
            $monitor("%b\t\t%b: %b",I, S, Y);
        #1  S = 3'bxxx;     I = 8'bxxxxxxxx;  

        #1  S = 3'b000;     I = 8'b00000000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b00000001;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b00000010;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b00000100;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b00001000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;        

        #1  S = 3'b000;     I = 8'b00010000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b00100000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b01000000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;

        #1  S = 3'b000;     I = 8'b10000000;        
        #1  S = 3'b001;      
        #1  S = 3'b010;      
        #1  S = 3'b011;      
        #1  S = 3'b100;      
        #1  S = 3'b101;      
        #1  S = 3'b110;      
        #1  S = 3'b111;
        #1  $stop;
        
    end
            


    
endmodule