module test;
    reg A, B, X, Y;

    initial begin
       $monitor("%0b %0b %0b %0b", A, B, C, D);
       
    end

endmodule;